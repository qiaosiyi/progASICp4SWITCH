`timescale 1ns / 1ps
//pkt_ctl 0x00:invalid
//pkt_ctl 0x01:start
//pkt_ctl 0x02:stop
//pkt_ctl 0x03:64byte packet, only takes one cycle.


module test_b;

	wire out_valid_pid;
	wire [8:0] out_pid;
	wire [511:0] header;
	
	reg	reset=1, clk=0;
	reg [511:0] pkt_data [0:49];
	reg [7:0] pkt_ctl [0:49];
	reg [0:0] times=0;
	reg [7:0] pkt_cnt=0;
	
	reg in_valid_pkt=0;
	reg [7:0] in_pkt_ctl=0;
	reg [511:0] in_pkt_data=0;
	
	
	always begin
		#5 clk = 1;
		#5 clk = 0;
	end

	initial begin

		#7 reset = 1;

		#23 reset = 0;
	end
   
   
always@(posedge clk or reset)begin
		if(reset)begin
			pkt_ctl[ 0 ] = 1 ; pkt_data[0] ='h645464e4548454f4540200000000000010000110e62e6dbca30098009800ff9261ca079261ca7c4311080000c3a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 1 ] = 3 ; pkt_data[1] ='h100002000014141434d4540554a4647454346484643464b454945434; pkt_ctl[ 2 ] = 1 ; pkt_data[2] ='h54e4547454545454540200000000000010000110a62e3efea30098009800ff9261ca079261ca6c4311080000d3a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 3 ] = 3 ; pkt_data[3] ='h100002000014141434143414341434b454846434541464a4648454e4; pkt_ctl[ 4 ] = 1 ; pkt_data[4] ='h649464a464545444540200000000000010000110962e0efda30098009800ff9261ca079261ca5c4311080000e3a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 5 ] = 3 ; pkt_data[5] ='h10000200001414143414341434d454c454e454d45444646454446494; pkt_ctl[ 6 ] = 1 ; pkt_data[6] ='h649464a464545444540200000000000010000110962e0efda30098009800ff9261ca079261caeb431108000054a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 7 ] = 3 ; pkt_data[7] ='h10000200001414143414341434d454c454e454d45444646454446494; pkt_ctl[ 8 ] = 1 ; pkt_data[8] ='h54e4547454545454540200000000000010000110a62e3efea30098009800ff9261ca079261cadb431108000064a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 9 ] = 3 ; pkt_data[9] ='h100002000014141434143414341434b454846434541464a4648454e4; pkt_ctl[ 10 ] = 1 ; pkt_data[10] ='h645464e4548454f4540200000000000010000110e62e6dbca30098009800ff9261ca079261cacb431108000074a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 11 ] = 3 ; pkt_data[11] ='h100002000014141434d4540554a4647454346484643464b454945434; pkt_ctl[ 12 ] = 1 ; pkt_data[12] ='h645464e4548454f4540200000000000010000110e62e6dbca30098009800ff9261ca079261ca1b431108000025a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 13 ] = 3 ; pkt_data[13] ='h100002000014141434d4540554a4647454346484643464b454945434; pkt_ctl[ 14 ] = 1 ; pkt_data[14] ='h54e4547454545454540200000000000010000110a62e3efea30098009800ff9261ca079261ca0b431108000035a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 15 ] = 3 ; pkt_data[15] ='h100002000014141434143414341434b454846434541464a4648454e4; pkt_ctl[ 16 ] = 1 ; pkt_data[16] ='h649464a464545444540200000000000010000110962e0efda30098009800ff9261ca079261cafa431108000045a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 17 ] = 3 ; pkt_data[17] ='h10000200001414143414341434d454c454e454d45444646454446494; pkt_ctl[ 18 ] = 4 ; pkt_data[18] ='h000000000000000000000000000000000000ef9261ca000000000000249261ca684b52e01f8210004060008010006080684b52e01f82ffffffffffff; pkt_ctl[ 19 ] = 1 ; pkt_data[19] ='h54546424544464a4540200000000000010000110272e6e82a30098009800ff9261ca079261ca9a4311080000a5a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 20 ] = 3 ; pkt_data[20] ='h10000200001414143414341434143414341434143414341434146424; pkt_ctl[ 21 ] = 1 ; pkt_data[21] ='h54546424544464a4540200000000000010000110272e6e82a30098009800ff9261ca079261ca8a4311080000b5a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 22 ] = 3 ; pkt_data[22] ='h10000200001414143414341434143414341434143414341434146424; pkt_ctl[ 23 ] = 4 ; pkt_data[23] ='h0000000000000000000000000000000000004a9261ca371dd8a79b4e000000004acfff3e8000100040600080100060804acfff3e8000371dd8a79b4e; pkt_ctl[ 24 ] = 4 ; pkt_data[24] ='h000000004acfff3e80004a9261ca371dd8a79b4e20004060008010006080371dd8a79b4e4acfff3e8000; pkt_ctl[ 25 ] = 4 ; pkt_data[25] ='h000000ee52ff7001051ddbab62ee28262709f1cd8d104a61ca4a9261ca0000600800049d91920000540080371dd8a79b4e09dfff3e8000; pkt_ctl[ 26 ] = 4 ; pkt_data[26] ='h00000000000000008af9f0810105fe2826271ddbab62cd8d09f14a9261ca104a61cad1b460c300001ed082000054008009dfff3e8000371dd8a79b4e; pkt_ctl[ 27 ] = 1 ; pkt_data[27] ='h54546424544464a4540200000000000010000110272e6e82a30098009800ff9261ca079261ca0a431108000036a5e400005400809e8354e01f82ffffffffffff; pkt_ctl[ 28 ] = 3 ; pkt_data[28] ='h10000200001414143414341434143414341434143414341434146424; pkt_ctl[ 29 ] = 4 ; pkt_data[29] ='h0000009681ff000105aeb48251c863dba17800938fc76961ca4a9261ca0000600800040950920000540080371dd8a79b4e09dfff3e8000; pkt_ctl[ 30 ] = 1 ; pkt_data[30] ='hdba1c863dba1a050101000000c21ff000108d863dba1aeb48251938f78004a9261cac76961ca1e3960d70004591543000054008009dfff3e8000371dd8a79b4e; pkt_ctl[ 31 ] = 3 ; pkt_data[31] ='hd863; pkt_ctl[ 32 ] = 4 ; pkt_data[32] ='h0000000000000000a6beff000105d863dba19eb48251938f78004a9261cac76961caae3960d70004791592000054008009dfff3e8000371dd8a79b4e; pkt_ctl[ 33 ] = 1 ; pkt_data[33] ='h82519eb48251a050101000004781ff000108aeb48251d863dba17800938fc76961ca4a9261ca0000600800041950430000540080371dd8a79b4e09dfff3e8000; pkt_ctl[ 34 ] = 3 ; pkt_data[34] ='haeb4; pkt_ctl[ 35 ] = 4 ; pkt_data[35] ='h0000000000000000d396001001052d489080cfe11d8ac38f260e4a9261cac76961ca4e3960d70004d91592000054008009dfff3e8000371dd8a79b4e; pkt_ctl[ 36 ] = 1 ; pkt_data[36] ='h1d8acfe11d8aa05010100000478120800108dfe11d8a2d489080260ec38fc76961ca4a9261ca0000600800042950430000540080371dd8a79b4e09dfff3e8000; pkt_ctl[ 37 ] = 3 ; pkt_data[37] ='hdfe1; pkt_ctl[ 38 ] = 4 ; pkt_data[38] ='h0000000000000000cbc2bf00010567e9b95689bb681da38f260e4a9261cac76961ca3e3960d70004e91592000054008009dfff3e8000371dd8a79b4e; pkt_ctl[ 39 ] = 1 ; pkt_data[39] ='h681d89bb681da0501010000047813080010899bb681d67e9b956260ea38fc76961ca4a9261ca0000600800043950430000540080371dd8a79b4e09dfff3e8000; pkt_ctl[ 40 ] = 3 ; pkt_data[40] ='h99bb; pkt_ctl[ 41 ] = 1 ; pkt_data[41] ='h000000000062003030710000086affff81053023f22f0f39d701be9cbb104a9261ca2ed1468235ed60f60004151135000054008009dfff3e8000371dd8a79b4e; pkt_ctl[ 42 ] = 3 ; pkt_data[42] ='hb10ebff3cf81d92d1b1588bff6271a02977e90c4cf0ee82b765f540f32b3d32000; pkt_ctl[ 43 ] = 1 ; pkt_data[43] ='h0000000000620030307100002fc7204081055e21f896304b5a96968dbb104a9261ca262426435a3a6007000418a135000054008009dfff3e8000371dd8a79b4e; pkt_ctl[ 44 ] = 3 ; pkt_data[44] ='h066a11ec09489ac65fd36404992b92394d0b40ba600c11f9df2b874cc1c8ef0000; pkt_ctl[ 45 ] = 1 ; pkt_data[45] ='h54146424549464020000bb00a800589261ca60bbe011ed9e1d00a800a800ff9261ca589261ca18e0110800006df75e00005400806dff512fbd81ffffffffffff; pkt_ctl[ 46 ] = 2 ; pkt_data[46] ='h24d435ff00e424143414341434143414341434143414341434143414349464f454d45494640200143414341434244444445454f4542454f4542454a464245454; pkt_ctl[ 47 ] = 2 ; pkt_data[47] ='h230020000000100030006500120000000000000000308e0000000000000000001200001100000000000000000000000000000000000000000000000000000052; pkt_ctl[ 48 ] = 3 ; pkt_data[48] ='h00aa5510f0001001301060000000133344e414e41495144405148500a0cf08001000543575f42524c545f4c435c49414d4c500; pkt_ctl[ 49 ] = 4 ; pkt_data[49] ='h0000b1c1ff000105b149d7013023f22fbb10be9c2ed146824a9261ca0000600800041c60820000540080371dd8a79b4e09dfff3e8000; pkt_ctl[ 50 ] = 4 ; pkt_data[50] ='h000099c4ef000105e24b5a965e21f896bb10968d262426434a9261ca0000600800047e27820000540080371dd8a79b4e09dfff3e8000;
		end else begin
			if(times == 1)begin
				in_pkt_data <= pkt_data[pkt_cnt];
				in_pkt_ctl <= pkt_ctl[pkt_cnt];
				in_valid_pkt <= 1;
				pkt_cnt <= pkt_cnt + 1;
			end else begin
				in_pkt_ctl <= 0;
				in_valid_pkt <= 0;
			end
			times <= times + 1;
		end
	end
	
	mmu #(
		
	) mmu_inst(
		.clk(clk),
		.reset(reset),
		.in_valid_pkt_fifo(in_valid_pkt),
		.in_pkt_ctl_fifo(in_pkt_ctl),
		.in_pkt_data_fifo(in_pkt_data),
		
		.in_valid_pid_fifo(),
		.in_pid_fifo(),
		.in_pid_valid_lenth_fifo(),//有效长度*512等于发送出去的长度。
		
		.out_valid_pid(out_valid_pid),
		.out_pid(out_pid),
		.header(header)
	);
	

endmodule // main
