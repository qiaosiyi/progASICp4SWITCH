`timescale 1ps/1ps
module mp{
input               flow_id_vld_in,
input               flow_id_is_rx_in,
input               flow_id_match_in,
input   [22:0]      flow_id_in,

input               tx_flow_state_in_VALID,
input   [31:0]      tx_flow_state_in_DATA,
input               rx_flow_state_in_VALID,
input   [64:0]      rx_flow_state_in_DATA,

};

endmodule
