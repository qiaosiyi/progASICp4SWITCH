`timescale 1ns / 1ps

module probability #(
  parameter  C_LENGTH_WIDTH = 16,
  parameter  C_ID_WIDTH = 12,
  parameter  C_COUNTER_WIDTH = 20,
  parameter  C_pd_WIDTH = 32
  )(
    
    
  input                                         in_next_valid,
  input                   [C_LENGTH_WIDTH-1:0]  in_next_length,     //packets lenth value
  input                       [C_ID_WIDTH-1:0]  in_next_id,       //packets FLOW-ID
  input                  [C_COUNTER_WIDTH-1:0]  in_next_counter,     //counter value for index ID
  
  input                                       in_set_plut_valid, //BRAM INTERFACE
  input                       [11:0]            in_set_pult_add,
  input                       [31:0]           in_set_pult_value,
  
  output reg                                    out_couter_update_valid,
  output reg             [C_COUNTER_WIDTH-1:0]  out_counter_data_new,
  output reg                                    out_pd_valid,
  output reg                  [C_pd_WIDTH-1:0]  out_pd_data,
  output reg                  [C_ID_WIDTH-1:0]  out_id_data_next,    //if any valid signals include 1,out_couter_update_valid 2,out_pd_valid. "out_id_data_next"should be valid too.
	
  input                                         clk,
  input                                         rst
  );
  
  reg                                   [23:0]  PLUT  [1250:3072];
  reg                                   [23:0]  pd_data_tmp;
  reg                     [C_LENGTH_WIDTH-1:0]  next_length_tmp;
  reg                                    [8:0]  pre_state;
  reg                                    [8:0]  next_state;
  
  reg                                          set_plut_down;
  reg                            [11:0]  lookup_add_bram;
  wire                           [23:0]  lookup_data_bram;
  
  localparam                                    S_IDLE = 0;
  localparam                                    S_ADD = 1;
  localparam                                    S_INITIAL = 2;
  localparam                                    S_CALCMUL = 3;
  localparam                                    S_RESET = 4;
  localparam                                    S_ENABLE = 5;
  localparam                                    S_LOOKUP = 6;
  localparam                                    S_CALCMUL2 = 7;
  localparam                                    C_MAGIC_NUMBER = 292738;
  
  blk_mem_gen_4096_24 bram_plut_inst(               
    .clka(clk),              
    .ena(in_set_plut_valid),              
    .wea(1),              
    .addra(in_set_pult_add),            
    .dina(in_set_pult_value),              
    .douta(),            
    .clkb(clk),                       
    .enb(1),         
    .web(0),         
    .addrb(lookup_add_bram),       
    .dinb(),         
    .doutb(lookup_data_bram)       
  );  
  always @(posedge clk)begin
      if(rst)begin
	      set_plut_down <= 0;
	  end else begin
	      if(in_set_plut_valid)begin
		      set_plut_down <= 1;
		  end
	  end
  end

//////////////===============================FSM1========================================
  always @ (posedge clk) begin
    if (rst) begin
      pre_state <= S_IDLE;
    end else begin
      pre_state <= next_state;
    end
  end  
//////////////================================FSM2=======================================
  always @ (*) begin
    case(pre_state)//pre_state
      S_IDLE: begin
        if(in_next_valid)begin
          if(in_next_counter < C_MAGIC_NUMBER )begin             //if counter value is a small number, counter should be line way adding
            next_state = S_ADD;
          end else if(in_next_counter < 20'b1000_0000_0000_0000_0000) begin    //if C_Data should be inited, 20bits = 1 + 19 bits
            next_state = S_INITIAL;
          end else if(set_plut_down == 0) begin                    //counter value is large number 
            next_state = S_CALCMUL;
          end else begin
		    next_state = S_ENABLE;
		  end
        end else begin
          next_state = S_IDLE;
        end
      end
      S_ADD: begin
        next_state = S_IDLE;
      end
      S_INITIAL: begin
        next_state = S_IDLE;
      end
      S_CALCMUL: begin
        next_state = S_RESET;
      end
	  S_ENABLE: begin
        next_state = S_LOOKUP;
      end
	  S_LOOKUP: begin
        next_state = S_CALCMUL2;
      end
	  S_CALCMUL2: begin
        next_state = S_RESET;
      end
      S_RESET: begin
        next_state = S_IDLE;
      end
    endcase
  end  

//////////////=============================FSM3==========================================

  always @(posedge clk ) begin
    if(rst)begin
      PLUT[1250] <= 2429315;PLUT[1251] <= 2414826;PLUT[1252] <= 2400424;PLUT[1253] <= 2386107;PLUT[1254] <= 2371876;PLUT[1255] <= 2357729;PLUT[1256] <= 2343667;PLUT[1257] <= 2329689;PLUT[1258] <= 2315795;PLUT[1259] <= 2301983;PLUT[1260] <= 2288253;PLUT[1261] <= 2274605;PLUT[1262] <= 2261039;PLUT[1263] <= 2247554;PLUT[1264] <= 2234149;PLUT[1265] <= 2220824;PLUT[1266] <= 2207579;PLUT[1267] <= 2194412;PLUT[1268] <= 2181324;PLUT[1269] <= 2168314;PLUT[1270] <= 2155382;PLUT[1271] <= 2142527;PLUT[1272] <= 2129748;PLUT[1273] <= 2117046;PLUT[1274] <= 2104420;PLUT[1275] <= 2091868;PLUT[1276] <= 2079392;PLUT[1277] <= 2066990;PLUT[1278] <= 2054662;PLUT[1279] <= 2042408;PLUT[1280] <= 2030226;PLUT[1281] <= 2018118;PLUT[1282] <= 2006081;PLUT[1283] <= 1994116;PLUT[1284] <= 1982223;PLUT[1285] <= 1970401;PLUT[1286] <= 1958649;PLUT[1287] <= 1946967;PLUT[1288] <= 1935355;PLUT[1289] <= 1923812;PLUT[1290] <= 1912338;PLUT[1291] <= 1900932;PLUT[1292] <= 1889595;PLUT[1293] <= 1878325;PLUT[1294] <= 1867122;PLUT[1295] <= 1855986;PLUT[1296] <= 1844917;PLUT[1297] <= 1833913;PLUT[1298] <= 1822975;PLUT[1299] <= 1812103;PLUT[1300] <= 1801295;PLUT[1301] <= 1790552;PLUT[1302] <= 1779872;PLUT[1303] <= 1769257;PLUT[1304] <= 1758705;PLUT[1305] <= 1748215;PLUT[1306] <= 1737788;PLUT[1307] <= 1727424;PLUT[1308] <= 1717121;PLUT[1309] <= 1706880;PLUT[1310] <= 1696700;PLUT[1311] <= 1686580;PLUT[1312] <= 1676521;PLUT[1313] <= 1666522;PLUT[1314] <= 1656582;PLUT[1315] <= 1646702;PLUT[1316] <= 1636881;PLUT[1317] <= 1627118;PLUT[1318] <= 1617414;PLUT[1319] <= 1607767;PLUT[1320] <= 1598178;PLUT[1321] <= 1588646;PLUT[1322] <= 1579171;PLUT[1323] <= 1569753;PLUT[1324] <= 1560390;PLUT[1325] <= 1551084;PLUT[1326] <= 1541833;PLUT[1327] <= 1532637;PLUT[1328] <= 1523496;PLUT[1329] <= 1514410;PLUT[1330] <= 1505377;PLUT[1331] <= 1496399;PLUT[1332] <= 1487474;PLUT[1333] <= 1478602;PLUT[1334] <= 1469784;PLUT[1335] <= 1461018;PLUT[1336] <= 1452304;PLUT[1337] <= 1443642;PLUT[1338] <= 1435032;PLUT[1339] <= 1426473;PLUT[1340] <= 1417965;PLUT[1341] <= 1409508;PLUT[1342] <= 1401101;PLUT[1343] <= 1392745;PLUT[1344] <= 1384438;PLUT[1345] <= 1376181;PLUT[1346] <= 1367973;PLUT[1347] <= 1359815;PLUT[1348] <= 1351704;PLUT[1349] <= 1343642;PLUT[1350] <= 1335629;PLUT[1351] <= 1327663;PLUT[1352] <= 1319744;PLUT[1353] <= 1311873;PLUT[1354] <= 1304049;PLUT[1355] <= 1296271;PLUT[1356] <= 1288540;PLUT[1357] <= 1280855;PLUT[1358] <= 1273215;PLUT[1359] <= 1265622;PLUT[1360] <= 1258073;PLUT[1361] <= 1250570;PLUT[1362] <= 1243111;PLUT[1363] <= 1235697;PLUT[1364] <= 1228327;PLUT[1365] <= 1221001;PLUT[1366] <= 1213719;PLUT[1367] <= 1206480;PLUT[1368] <= 1199284;PLUT[1369] <= 1192131;PLUT[1370] <= 1185021;PLUT[1371] <= 1177953;PLUT[1372] <= 1170928;PLUT[1373] <= 1163944;PLUT[1374] <= 1157002;PLUT[1375] <= 1150102;PLUT[1376] <= 1143242;PLUT[1377] <= 1136424;PLUT[1378] <= 1129646;PLUT[1379] <= 1122908;PLUT[1380] <= 1116211;PLUT[1381] <= 1109554;PLUT[1382] <= 1102936;PLUT[1383] <= 1096358;PLUT[1384] <= 1089819;PLUT[1385] <= 1083319;PLUT[1386] <= 1076858;PLUT[1387] <= 1070435;PLUT[1388] <= 1064051;PLUT[1389] <= 1057705;PLUT[1390] <= 1051396;PLUT[1391] <= 1045126;PLUT[1392] <= 1038892;PLUT[1393] <= 1032696;PLUT[1394] <= 1026537;PLUT[1395] <= 1020414;PLUT[1396] <= 1014328;PLUT[1397] <= 1008279;PLUT[1398] <= 1002265;PLUT[1399] <= 996287;PLUT[1400] <= 990345;PLUT[1401] <= 984439;PLUT[1402] <= 978567;PLUT[1403] <= 972731;PLUT[1404] <= 966929;PLUT[1405] <= 961162;PLUT[1406] <= 955430;PLUT[1407] <= 949731;PLUT[1408] <= 944067;PLUT[1409] <= 938436;PLUT[1410] <= 932839;PLUT[1411] <= 927276;PLUT[1412] <= 921745;PLUT[1413] <= 916248;PLUT[1414] <= 910783;PLUT[1415] <= 905351;PLUT[1416] <= 899951;PLUT[1417] <= 894584;PLUT[1418] <= 889248;PLUT[1419] <= 883944;PLUT[1420] <= 878672;PLUT[1421] <= 873432;PLUT[1422] <= 868222;PLUT[1423] <= 863044;PLUT[1424] <= 857897;PLUT[1425] <= 852780;PLUT[1426] <= 847694;PLUT[1427] <= 842638;PLUT[1428] <= 837612;PLUT[1429] <= 832617;PLUT[1430] <= 827651;PLUT[1431] <= 822715;PLUT[1432] <= 817808;PLUT[1433] <= 812930;PLUT[1434] <= 808082;PLUT[1435] <= 803262;PLUT[1436] <= 798471;PLUT[1437] <= 793709;PLUT[1438] <= 788975;PLUT[1439] <= 784270;PLUT[1440] <= 779592;PLUT[1441] <= 774942;PLUT[1442] <= 770320;PLUT[1443] <= 765726;PLUT[1444] <= 761159;PLUT[1445] <= 756619;PLUT[1446] <= 752107;PLUT[1447] <= 747621;PLUT[1448] <= 743162;PLUT[1449] <= 738730;PLUT[1450] <= 734324;PLUT[1451] <= 729944;PLUT[1452] <= 725590;PLUT[1453] <= 721263;PLUT[1454] <= 716961;PLUT[1455] <= 712685;PLUT[1456] <= 708434;PLUT[1457] <= 704209;PLUT[1458] <= 700009;PLUT[1459] <= 695834;PLUT[1460] <= 691684;PLUT[1461] <= 687559;PLUT[1462] <= 683458;PLUT[1463] <= 679382;PLUT[1464] <= 675330;PLUT[1465] <= 671302;PLUT[1466] <= 667298;PLUT[1467] <= 663318;PLUT[1468] <= 659362;PLUT[1469] <= 655429;PLUT[1470] <= 651520;PLUT[1471] <= 647634;PLUT[1472] <= 643772;PLUT[1473] <= 639932;PLUT[1474] <= 636115;PLUT[1475] <= 632322;PLUT[1476] <= 628550;PLUT[1477] <= 624801;PLUT[1478] <= 621075;PLUT[1479] <= 617371;PLUT[1480] <= 613689;PLUT[1481] <= 610028;PLUT[1482] <= 606390;PLUT[1483] <= 602773;PLUT[1484] <= 599178;PLUT[1485] <= 595605;PLUT[1486] <= 592052;PLUT[1487] <= 588521;PLUT[1488] <= 585011;PLUT[1489] <= 581522;PLUT[1490] <= 578054;PLUT[1491] <= 574606;PLUT[1492] <= 571179;PLUT[1493] <= 567772;PLUT[1494] <= 564386;PLUT[1495] <= 561020;PLUT[1496] <= 557674;PLUT[1497] <= 554348;PLUT[1498] <= 551042;PLUT[1499] <= 547755;PLUT[1500] <= 544488;PLUT[1501] <= 541241;PLUT[1502] <= 538013;PLUT[1503] <= 534804;PLUT[1504] <= 531614;PLUT[1505] <= 528443;PLUT[1506] <= 525292;PLUT[1507] <= 522159;PLUT[1508] <= 519044;PLUT[1509] <= 515949;PLUT[1510] <= 512871;PLUT[1511] <= 509813;PLUT[1512] <= 506772;PLUT[1513] <= 503749;PLUT[1514] <= 500745;PLUT[1515] <= 497758;PLUT[1516] <= 494790;PLUT[1517] <= 491839;PLUT[1518] <= 488905;PLUT[1519] <= 485989;PLUT[1520] <= 483091;PLUT[1521] <= 480209;PLUT[1522] <= 477345;PLUT[1523] <= 474498;PLUT[1524] <= 471668;PLUT[1525] <= 468855;PLUT[1526] <= 466059;PLUT[1527] <= 463279;PLUT[1528] <= 460516;PLUT[1529] <= 457770;PLUT[1530] <= 455039;PLUT[1531] <= 452325;PLUT[1532] <= 449628;PLUT[1533] <= 446946;PLUT[1534] <= 444280;PLUT[1535] <= 441630;PLUT[1536] <= 438996;PLUT[1537] <= 436378;PLUT[1538] <= 433775;PLUT[1539] <= 431188;PLUT[1540] <= 428617;PLUT[1541] <= 426060;PLUT[1542] <= 423519;PLUT[1543] <= 420993;PLUT[1544] <= 418482;PLUT[1545] <= 415986;PLUT[1546] <= 413505;PLUT[1547] <= 411039;PLUT[1548] <= 408588;PLUT[1549] <= 406151;PLUT[1550] <= 403728;PLUT[1551] <= 401320;PLUT[1552] <= 398927;PLUT[1553] <= 396548;PLUT[1554] <= 394182;PLUT[1555] <= 391831;PLUT[1556] <= 389494;PLUT[1557] <= 387171;PLUT[1558] <= 384862;PLUT[1559] <= 382567;PLUT[1560] <= 380285;PLUT[1561] <= 378017;PLUT[1562] <= 375762;PLUT[1563] <= 373521;PLUT[1564] <= 371294;PLUT[1565] <= 369079;PLUT[1566] <= 366878;PLUT[1567] <= 364690;PLUT[1568] <= 362515;PLUT[1569] <= 360352;PLUT[1570] <= 358203;PLUT[1571] <= 356067;PLUT[1572] <= 353943;PLUT[1573] <= 351832;PLUT[1574] <= 349734;PLUT[1575] <= 347648;PLUT[1576] <= 345574;PLUT[1577] <= 343513;PLUT[1578] <= 341465;PLUT[1579] <= 339428;PLUT[1580] <= 337404;PLUT[1581] <= 335391;PLUT[1582] <= 333391;PLUT[1583] <= 331402;PLUT[1584] <= 329426;PLUT[1585] <= 327461;PLUT[1586] <= 325508;PLUT[1587] <= 323567;PLUT[1588] <= 321637;PLUT[1589] <= 319719;PLUT[1590] <= 317812;PLUT[1591] <= 315916;PLUT[1592] <= 314032;PLUT[1593] <= 312159;PLUT[1594] <= 310297;PLUT[1595] <= 308447;PLUT[1596] <= 306607;PLUT[1597] <= 304778;PLUT[1598] <= 302960;PLUT[1599] <= 301154;PLUT[1600] <= 299357;PLUT[1601] <= 297572;PLUT[1602] <= 295797;PLUT[1603] <= 294033;PLUT[1604] <= 292279;PLUT[1605] <= 290536;PLUT[1606] <= 288803;PLUT[1607] <= 287081;PLUT[1608] <= 285369;PLUT[1609] <= 283667;PLUT[1610] <= 281975;PLUT[1611] <= 280293;PLUT[1612] <= 278621;PLUT[1613] <= 276959;PLUT[1614] <= 275308;PLUT[1615] <= 273666;PLUT[1616] <= 272033;PLUT[1617] <= 270411;PLUT[1618] <= 268798;PLUT[1619] <= 267195;PLUT[1620] <= 265601;PLUT[1621] <= 264017;PLUT[1622] <= 262443;PLUT[1623] <= 260877;PLUT[1624] <= 259321;PLUT[1625] <= 257775;PLUT[1626] <= 256237;PLUT[1627] <= 254709;PLUT[1628] <= 253190;PLUT[1629] <= 251680;PLUT[1630] <= 250179;PLUT[1631] <= 248687;PLUT[1632] <= 247203;PLUT[1633] <= 245729;PLUT[1634] <= 244263;PLUT[1635] <= 242807;PLUT[1636] <= 241358;PLUT[1637] <= 239919;PLUT[1638] <= 238488;PLUT[1639] <= 237066;PLUT[1640] <= 235652;PLUT[1641] <= 234246;PLUT[1642] <= 232849;PLUT[1643] <= 231460;PLUT[1644] <= 230080;PLUT[1645] <= 228708;PLUT[1646] <= 227344;PLUT[1647] <= 225988;PLUT[1648] <= 224640;PLUT[1649] <= 223300;PLUT[1650] <= 221968;PLUT[1651] <= 220644;PLUT[1652] <= 219328;PLUT[1653] <= 218020;PLUT[1654] <= 216720;PLUT[1655] <= 215427;PLUT[1656] <= 214142;PLUT[1657] <= 212865;PLUT[1658] <= 211596;PLUT[1659] <= 210334;PLUT[1660] <= 209079;PLUT[1661] <= 207832;PLUT[1662] <= 206593;PLUT[1663] <= 205360;PLUT[1664] <= 204136;PLUT[1665] <= 202918;PLUT[1666] <= 201708;PLUT[1667] <= 200505;PLUT[1668] <= 199309;PLUT[1669] <= 198120;PLUT[1670] <= 196939;PLUT[1671] <= 195764;PLUT[1672] <= 194596;PLUT[1673] <= 193436;PLUT[1674] <= 192282;PLUT[1675] <= 191135;PLUT[1676] <= 189995;PLUT[1677] <= 188862;PLUT[1678] <= 187736;PLUT[1679] <= 186616;PLUT[1680] <= 185503;PLUT[1681] <= 184397;PLUT[1682] <= 183297;PLUT[1683] <= 182204;PLUT[1684] <= 181117;PLUT[1685] <= 180037;PLUT[1686] <= 178963;PLUT[1687] <= 177896;PLUT[1688] <= 176835;PLUT[1689] <= 175780;PLUT[1690] <= 174731;PLUT[1691] <= 173689;PLUT[1692] <= 172653;PLUT[1693] <= 171624;PLUT[1694] <= 170600;PLUT[1695] <= 169583;PLUT[1696] <= 168571;PLUT[1697] <= 167566;PLUT[1698] <= 166566;PLUT[1699] <= 165573;PLUT[1700] <= 164585;PLUT[1701] <= 163604;PLUT[1702] <= 162628;PLUT[1703] <= 161658;PLUT[1704] <= 160694;PLUT[1705] <= 159735;PLUT[1706] <= 158783;PLUT[1707] <= 157836;PLUT[1708] <= 156894;PLUT[1709] <= 155959;PLUT[1710] <= 155028;PLUT[1711] <= 154104;PLUT[1712] <= 153185;PLUT[1713] <= 152271;PLUT[1714] <= 151363;PLUT[1715] <= 150460;PLUT[1716] <= 149563;PLUT[1717] <= 148671;PLUT[1718] <= 147784;PLUT[1719] <= 146903;PLUT[1720] <= 146026;PLUT[1721] <= 145156;PLUT[1722] <= 144290;PLUT[1723] <= 143429;PLUT[1724] <= 142574;PLUT[1725] <= 141723;PLUT[1726] <= 140878;PLUT[1727] <= 140038;PLUT[1728] <= 139203;PLUT[1729] <= 138372;PLUT[1730] <= 137547;PLUT[1731] <= 136727;PLUT[1732] <= 135911;PLUT[1733] <= 135101;PLUT[1734] <= 134295;PLUT[1735] <= 133494;PLUT[1736] <= 132698;PLUT[1737] <= 131906;PLUT[1738] <= 131120;PLUT[1739] <= 130338;PLUT[1740] <= 129560;PLUT[1741] <= 128788;PLUT[1742] <= 128019;PLUT[1743] <= 127256;PLUT[1744] <= 126497;PLUT[1745] <= 125742;PLUT[1746] <= 124992;PLUT[1747] <= 124247;PLUT[1748] <= 123506;PLUT[1749] <= 122769;PLUT[1750] <= 122037;PLUT[1751] <= 121309;PLUT[1752] <= 120586;PLUT[1753] <= 119867;PLUT[1754] <= 119152;PLUT[1755] <= 118441;PLUT[1756] <= 117735;PLUT[1757] <= 117032;PLUT[1758] <= 116334;PLUT[1759] <= 115640;PLUT[1760] <= 114951;PLUT[1761] <= 114265;PLUT[1762] <= 113584;PLUT[1763] <= 112906;PLUT[1764] <= 112233;PLUT[1765] <= 111563;PLUT[1766] <= 110898;PLUT[1767] <= 110237;PLUT[1768] <= 109579;PLUT[1769] <= 108926;PLUT[1770] <= 108276;PLUT[1771] <= 107630;PLUT[1772] <= 106988;PLUT[1773] <= 106350;PLUT[1774] <= 105716;PLUT[1775] <= 105085;PLUT[1776] <= 104459;PLUT[1777] <= 103836;PLUT[1778] <= 103216;PLUT[1779] <= 102601;PLUT[1780] <= 101989;PLUT[1781] <= 101380;PLUT[1782] <= 100776;PLUT[1783] <= 100175;PLUT[1784] <= 99577;PLUT[1785] <= 98983;PLUT[1786] <= 98393;PLUT[1787] <= 97806;PLUT[1788] <= 97223;PLUT[1789] <= 96643;PLUT[1790] <= 96067;PLUT[1791] <= 95494;PLUT[1792] <= 94924;PLUT[1793] <= 94358;PLUT[1794] <= 93795;PLUT[1795] <= 93236;PLUT[1796] <= 92680;PLUT[1797] <= 92127;PLUT[1798] <= 91577;PLUT[1799] <= 91031;PLUT[1800] <= 90488;PLUT[1801] <= 89949;PLUT[1802] <= 89412;PLUT[1803] <= 88879;PLUT[1804] <= 88349;PLUT[1805] <= 87822;PLUT[1806] <= 87298;PLUT[1807] <= 86777;PLUT[1808] <= 86260;PLUT[1809] <= 85745;PLUT[1810] <= 85234;PLUT[1811] <= 84726;PLUT[1812] <= 84220;PLUT[1813] <= 83718;PLUT[1814] <= 83219;PLUT[1815] <= 82722;PLUT[1816] <= 82229;PLUT[1817] <= 81738;PLUT[1818] <= 81251;PLUT[1819] <= 80766;PLUT[1820] <= 80285;PLUT[1821] <= 79806;PLUT[1822] <= 79330;PLUT[1823] <= 78857;PLUT[1824] <= 78386;PLUT[1825] <= 77919;PLUT[1826] <= 77454;PLUT[1827] <= 76992;PLUT[1828] <= 76533;PLUT[1829] <= 76076;PLUT[1830] <= 75623;PLUT[1831] <= 75172;PLUT[1832] <= 74723;PLUT[1833] <= 74278;PLUT[1834] <= 73835;PLUT[1835] <= 73394;PLUT[1836] <= 72957;PLUT[1837] <= 72521;PLUT[1838] <= 72089;PLUT[1839] <= 71659;PLUT[1840] <= 71232;PLUT[1841] <= 70807;PLUT[1842] <= 70384;PLUT[1843] <= 69965;PLUT[1844] <= 69547;PLUT[1845] <= 69133;PLUT[1846] <= 68720;PLUT[1847] <= 68310;PLUT[1848] <= 67903;PLUT[1849] <= 67498;PLUT[1850] <= 67095;PLUT[1851] <= 66695;PLUT[1852] <= 66297;PLUT[1853] <= 65902;PLUT[1854] <= 65509;PLUT[1855] <= 65118;PLUT[1856] <= 64730;PLUT[1857] <= 64344;PLUT[1858] <= 63960;PLUT[1859] <= 63579;PLUT[1860] <= 63199;PLUT[1861] <= 62822;PLUT[1862] <= 62448;PLUT[1863] <= 62075;PLUT[1864] <= 61705;PLUT[1865] <= 61337;PLUT[1866] <= 60971;PLUT[1867] <= 60607;PLUT[1868] <= 60246;PLUT[1869] <= 59887;PLUT[1870] <= 59530;PLUT[1871] <= 59174;PLUT[1872] <= 58822;PLUT[1873] <= 58471;PLUT[1874] <= 58122;PLUT[1875] <= 57775;PLUT[1876] <= 57431;PLUT[1877] <= 57088;PLUT[1878] <= 56748;PLUT[1879] <= 56409;PLUT[1880] <= 56073;PLUT[1881] <= 55738;PLUT[1882] <= 55406;PLUT[1883] <= 55075;PLUT[1884] <= 54747;PLUT[1885] <= 54420;PLUT[1886] <= 54096;PLUT[1887] <= 53773;PLUT[1888] <= 53453;PLUT[1889] <= 53134;PLUT[1890] <= 52817;PLUT[1891] <= 52502;PLUT[1892] <= 52189;PLUT[1893] <= 51877;PLUT[1894] <= 51568;PLUT[1895] <= 51260;PLUT[1896] <= 50955;PLUT[1897] <= 50651;PLUT[1898] <= 50349;PLUT[1899] <= 50048;PLUT[1900] <= 49750;PLUT[1901] <= 49453;PLUT[1902] <= 49158;PLUT[1903] <= 48865;PLUT[1904] <= 48574;PLUT[1905] <= 48284;PLUT[1906] <= 47996;PLUT[1907] <= 47710;PLUT[1908] <= 47425;PLUT[1909] <= 47142;PLUT[1910] <= 46861;PLUT[1911] <= 46582;PLUT[1912] <= 46304;PLUT[1913] <= 46028;PLUT[1914] <= 45753;PLUT[1915] <= 45480;PLUT[1916] <= 45209;PLUT[1917] <= 44939;PLUT[1918] <= 44671;PLUT[1919] <= 44405;PLUT[1920] <= 44140;PLUT[1921] <= 43877;PLUT[1922] <= 43615;PLUT[1923] <= 43355;PLUT[1924] <= 43096;PLUT[1925] <= 42839;PLUT[1926] <= 42584;PLUT[1927] <= 42330;PLUT[1928] <= 42077;PLUT[1929] <= 41826;PLUT[1930] <= 41577;PLUT[1931] <= 41329;PLUT[1932] <= 41082;PLUT[1933] <= 40837;PLUT[1934] <= 40594;PLUT[1935] <= 40352;PLUT[1936] <= 40111;PLUT[1937] <= 39872;PLUT[1938] <= 39634;PLUT[1939] <= 39398;PLUT[1940] <= 39163;PLUT[1941] <= 38929;PLUT[1942] <= 38697;PLUT[1943] <= 38466;PLUT[1944] <= 38237;PLUT[1945] <= 38009;PLUT[1946] <= 37782;PLUT[1947] <= 37557;PLUT[1948] <= 37333;PLUT[1949] <= 37110;PLUT[1950] <= 36889;PLUT[1951] <= 36669;PLUT[1952] <= 36450;PLUT[1953] <= 36232;PLUT[1954] <= 36016;PLUT[1955] <= 35802;PLUT[1956] <= 35588;PLUT[1957] <= 35376;PLUT[1958] <= 35165;PLUT[1959] <= 34955;PLUT[1960] <= 34747;PLUT[1961] <= 34539;PLUT[1962] <= 34333;PLUT[1963] <= 34129;PLUT[1964] <= 33925;PLUT[1965] <= 33723;PLUT[1966] <= 33521;PLUT[1967] <= 33322;PLUT[1968] <= 33123;PLUT[1969] <= 32925;PLUT[1970] <= 32729;PLUT[1971] <= 32534;PLUT[1972] <= 32340;PLUT[1973] <= 32147;PLUT[1974] <= 31955;PLUT[1975] <= 31764;PLUT[1976] <= 31575;PLUT[1977] <= 31387;PLUT[1978] <= 31199;PLUT[1979] <= 31013;PLUT[1980] <= 30828;PLUT[1981] <= 30645;PLUT[1982] <= 30462;PLUT[1983] <= 30280;PLUT[1984] <= 30099;PLUT[1985] <= 29920;PLUT[1986] <= 29741;PLUT[1987] <= 29564;PLUT[1988] <= 29388;PLUT[1989] <= 29213;PLUT[1990] <= 29038;PLUT[1991] <= 28865;PLUT[1992] <= 28693;PLUT[1993] <= 28522;PLUT[1994] <= 28352;PLUT[1995] <= 28183;PLUT[1996] <= 28014;PLUT[1997] <= 27847;PLUT[1998] <= 27681;PLUT[1999] <= 27516;PLUT[2000] <= 27352;PLUT[2001] <= 27189;PLUT[2002] <= 27027;PLUT[2003] <= 26866;PLUT[2004] <= 26705;PLUT[2005] <= 26546;PLUT[2006] <= 26388;PLUT[2007] <= 26230;PLUT[2008] <= 26074;PLUT[2009] <= 25918;PLUT[2010] <= 25764;PLUT[2011] <= 25610;PLUT[2012] <= 25457;PLUT[2013] <= 25306;PLUT[2014] <= 25155;PLUT[2015] <= 25005;PLUT[2016] <= 24855;PLUT[2017] <= 24707;PLUT[2018] <= 24560;PLUT[2019] <= 24413;PLUT[2020] <= 24268;PLUT[2021] <= 24123;PLUT[2022] <= 23979;PLUT[2023] <= 23836;PLUT[2024] <= 23694;PLUT[2025] <= 23553;PLUT[2026] <= 23412;PLUT[2027] <= 23273;PLUT[2028] <= 23134;PLUT[2029] <= 22996;PLUT[2030] <= 22859;PLUT[2031] <= 22722;PLUT[2032] <= 22587;PLUT[2033] <= 22452;PLUT[2034] <= 22318;PLUT[2035] <= 22185;PLUT[2036] <= 22053;PLUT[2037] <= 21921;PLUT[2038] <= 21790;PLUT[2039] <= 21660;PLUT[2040] <= 21531;PLUT[2041] <= 21403;PLUT[2042] <= 21275;PLUT[2043] <= 21148;PLUT[2044] <= 21022;PLUT[2045] <= 20897;PLUT[2046] <= 20772;PLUT[2047] <= 20648;PLUT[2048] <= 20525;PLUT[2049] <= 20403;PLUT[2050] <= 20281;PLUT[2051] <= 20160;PLUT[2052] <= 20040;PLUT[2053] <= 19920;PLUT[2054] <= 19801;PLUT[2055] <= 19683;PLUT[2056] <= 19566;PLUT[2057] <= 19449;PLUT[2058] <= 19333;PLUT[2059] <= 19218;PLUT[2060] <= 19103;PLUT[2061] <= 18989;PLUT[2062] <= 18876;PLUT[2063] <= 18764;PLUT[2064] <= 18652;PLUT[2065] <= 18540;PLUT[2066] <= 18430;PLUT[2067] <= 18320;PLUT[2068] <= 18211;PLUT[2069] <= 18102;PLUT[2070] <= 17994;PLUT[2071] <= 17887;PLUT[2072] <= 17780;PLUT[2073] <= 17674;PLUT[2074] <= 17569;PLUT[2075] <= 17464;PLUT[2076] <= 17360;PLUT[2077] <= 17256;PLUT[2078] <= 17153;PLUT[2079] <= 17051;PLUT[2080] <= 16949;PLUT[2081] <= 16848;PLUT[2082] <= 16748;PLUT[2083] <= 16648;PLUT[2084] <= 16548;PLUT[2085] <= 16450;PLUT[2086] <= 16352;PLUT[2087] <= 16254;PLUT[2088] <= 16157;PLUT[2089] <= 16061;PLUT[2090] <= 15965;PLUT[2091] <= 15870;PLUT[2092] <= 15775;PLUT[2093] <= 15681;PLUT[2094] <= 15587;PLUT[2095] <= 15494;PLUT[2096] <= 15402;PLUT[2097] <= 15310;PLUT[2098] <= 15219;PLUT[2099] <= 15128;PLUT[2100] <= 15038;PLUT[2101] <= 14948;PLUT[2102] <= 14859;PLUT[2103] <= 14770;PLUT[2104] <= 14682;PLUT[2105] <= 14595;PLUT[2106] <= 14508;PLUT[2107] <= 14421;PLUT[2108] <= 14335;PLUT[2109] <= 14250;PLUT[2110] <= 14165;PLUT[2111] <= 14080;PLUT[2112] <= 13996;PLUT[2113] <= 13913;PLUT[2114] <= 13830;PLUT[2115] <= 13747;PLUT[2116] <= 13665;PLUT[2117] <= 13584;PLUT[2118] <= 13503;PLUT[2119] <= 13422;PLUT[2120] <= 13342;PLUT[2121] <= 13263;PLUT[2122] <= 13183;PLUT[2123] <= 13105;PLUT[2124] <= 13027;PLUT[2125] <= 12949;PLUT[2126] <= 12872;PLUT[2127] <= 12795;PLUT[2128] <= 12719;PLUT[2129] <= 12643;PLUT[2130] <= 12567;PLUT[2131] <= 12492;PLUT[2132] <= 12418;PLUT[2133] <= 12344;PLUT[2134] <= 12270;PLUT[2135] <= 12197;PLUT[2136] <= 12124;PLUT[2137] <= 12052;PLUT[2138] <= 11980;PLUT[2139] <= 11909;PLUT[2140] <= 11838;PLUT[2141] <= 11767;PLUT[2142] <= 11697;PLUT[2143] <= 11627;PLUT[2144] <= 11558;PLUT[2145] <= 11489;PLUT[2146] <= 11420;PLUT[2147] <= 11352;PLUT[2148] <= 11284;PLUT[2149] <= 11217;PLUT[2150] <= 11150;PLUT[2151] <= 11084;PLUT[2152] <= 11018;PLUT[2153] <= 10952;PLUT[2154] <= 10887;PLUT[2155] <= 10822;PLUT[2156] <= 10757;PLUT[2157] <= 10693;PLUT[2158] <= 10629;PLUT[2159] <= 10566;PLUT[2160] <= 10503;PLUT[2161] <= 10440;PLUT[2162] <= 10378;PLUT[2163] <= 10316;PLUT[2164] <= 10254;PLUT[2165] <= 10193;PLUT[2166] <= 10132;PLUT[2167] <= 10072;PLUT[2168] <= 10012;PLUT[2169] <= 9952;PLUT[2170] <= 9893;PLUT[2171] <= 9834;PLUT[2172] <= 9775;PLUT[2173] <= 9717;PLUT[2174] <= 9659;PLUT[2175] <= 9601;PLUT[2176] <= 9544;PLUT[2177] <= 9487;PLUT[2178] <= 9431;PLUT[2179] <= 9374;PLUT[2180] <= 9318;PLUT[2181] <= 9263;PLUT[2182] <= 9208;PLUT[2183] <= 9153;PLUT[2184] <= 9098;PLUT[2185] <= 9044;PLUT[2186] <= 8990;PLUT[2187] <= 8936;PLUT[2188] <= 8883;PLUT[2189] <= 8830;PLUT[2190] <= 8777;PLUT[2191] <= 8725;PLUT[2192] <= 8673;PLUT[2193] <= 8621;PLUT[2194] <= 8570;PLUT[2195] <= 8519;PLUT[2196] <= 8468;PLUT[2197] <= 8417;PLUT[2198] <= 8367;PLUT[2199] <= 8317;PLUT[2200] <= 8268;PLUT[2201] <= 8218;PLUT[2202] <= 8169;PLUT[2203] <= 8120;PLUT[2204] <= 8072;PLUT[2205] <= 8024;PLUT[2206] <= 7976;PLUT[2207] <= 7928;PLUT[2208] <= 7881;PLUT[2209] <= 7834;PLUT[2210] <= 7787;PLUT[2211] <= 7741;PLUT[2212] <= 7695;PLUT[2213] <= 7649;PLUT[2214] <= 7603;PLUT[2215] <= 7558;PLUT[2216] <= 7513;PLUT[2217] <= 7468;PLUT[2218] <= 7424;PLUT[2219] <= 7379;PLUT[2220] <= 7335;PLUT[2221] <= 7291;PLUT[2222] <= 7248;PLUT[2223] <= 7205;PLUT[2224] <= 7162;PLUT[2225] <= 7119;PLUT[2226] <= 7077;PLUT[2227] <= 7034;PLUT[2228] <= 6992;PLUT[2229] <= 6951;PLUT[2230] <= 6909;PLUT[2231] <= 6868;PLUT[2232] <= 6827;PLUT[2233] <= 6786;PLUT[2234] <= 6746;PLUT[2235] <= 6706;PLUT[2236] <= 6666;PLUT[2237] <= 6626;PLUT[2238] <= 6586;PLUT[2239] <= 6547;PLUT[2240] <= 6508;PLUT[2241] <= 6469;PLUT[2242] <= 6431;PLUT[2243] <= 6392;PLUT[2244] <= 6354;PLUT[2245] <= 6316;PLUT[2246] <= 6279;PLUT[2247] <= 6241;PLUT[2248] <= 6204;PLUT[2249] <= 6167;PLUT[2250] <= 6130;PLUT[2251] <= 6094;PLUT[2252] <= 6057;PLUT[2253] <= 6021;PLUT[2254] <= 5985;PLUT[2255] <= 5949;PLUT[2256] <= 5914;PLUT[2257] <= 5879;PLUT[2258] <= 5844;PLUT[2259] <= 5809;PLUT[2260] <= 5774;PLUT[2261] <= 5740;PLUT[2262] <= 5705;PLUT[2263] <= 5671;PLUT[2264] <= 5638;PLUT[2265] <= 5604;PLUT[2266] <= 5571;PLUT[2267] <= 5537;PLUT[2268] <= 5504;PLUT[2269] <= 5471;PLUT[2270] <= 5439;PLUT[2271] <= 5406;PLUT[2272] <= 5374;PLUT[2273] <= 5342;PLUT[2274] <= 5310;PLUT[2275] <= 5279;PLUT[2276] <= 5247;PLUT[2277] <= 5216;PLUT[2278] <= 5185;PLUT[2279] <= 5154;PLUT[2280] <= 5123;PLUT[2281] <= 5092;PLUT[2282] <= 5062;PLUT[2283] <= 5032;PLUT[2284] <= 5002;PLUT[2285] <= 4972;PLUT[2286] <= 4942;PLUT[2287] <= 4913;PLUT[2288] <= 4884;PLUT[2289] <= 4854;PLUT[2290] <= 4825;PLUT[2291] <= 4797;PLUT[2292] <= 4768;PLUT[2293] <= 4740;PLUT[2294] <= 4711;PLUT[2295] <= 4683;PLUT[2296] <= 4655;PLUT[2297] <= 4628;PLUT[2298] <= 4600;PLUT[2299] <= 4573;PLUT[2300] <= 4545;PLUT[2301] <= 4518;PLUT[2302] <= 4491;PLUT[2303] <= 4464;PLUT[2304] <= 4438;PLUT[2305] <= 4411;PLUT[2306] <= 4385;PLUT[2307] <= 4359;PLUT[2308] <= 4333;PLUT[2309] <= 4307;PLUT[2310] <= 4281;PLUT[2311] <= 4256;PLUT[2312] <= 4230;PLUT[2313] <= 4205;PLUT[2314] <= 4180;PLUT[2315] <= 4155;PLUT[2316] <= 4130;PLUT[2317] <= 4106;PLUT[2318] <= 4081;PLUT[2319] <= 4057;PLUT[2320] <= 4033;PLUT[2321] <= 4009;PLUT[2322] <= 3985;PLUT[2323] <= 3961;PLUT[2324] <= 3937;PLUT[2325] <= 3914;PLUT[2326] <= 3890;PLUT[2327] <= 3867;PLUT[2328] <= 3844;PLUT[2329] <= 3821;PLUT[2330] <= 3798;PLUT[2331] <= 3776;PLUT[2332] <= 3753;PLUT[2333] <= 3731;PLUT[2334] <= 3709;PLUT[2335] <= 3687;PLUT[2336] <= 3665;PLUT[2337] <= 3643;PLUT[2338] <= 3621;PLUT[2339] <= 3599;PLUT[2340] <= 3578;PLUT[2341] <= 3557;PLUT[2342] <= 3535;PLUT[2343] <= 3514;PLUT[2344] <= 3493;PLUT[2345] <= 3472;PLUT[2346] <= 3452;PLUT[2347] <= 3431;PLUT[2348] <= 3411;PLUT[2349] <= 3390;PLUT[2350] <= 3370;PLUT[2351] <= 3350;PLUT[2352] <= 3330;PLUT[2353] <= 3310;PLUT[2354] <= 3290;PLUT[2355] <= 3271;PLUT[2356] <= 3251;PLUT[2357] <= 3232;PLUT[2358] <= 3213;PLUT[2359] <= 3193;PLUT[2360] <= 3174;PLUT[2361] <= 3155;PLUT[2362] <= 3137;PLUT[2363] <= 3118;PLUT[2364] <= 3099;PLUT[2365] <= 3081;PLUT[2366] <= 3062;PLUT[2367] <= 3044;PLUT[2368] <= 3026;PLUT[2369] <= 3008;PLUT[2370] <= 2990;PLUT[2371] <= 2972;PLUT[2372] <= 2954;PLUT[2373] <= 2937;PLUT[2374] <= 2919;PLUT[2375] <= 2902;PLUT[2376] <= 2885;PLUT[2377] <= 2867;PLUT[2378] <= 2850;PLUT[2379] <= 2833;PLUT[2380] <= 2816;PLUT[2381] <= 2800;PLUT[2382] <= 2783;PLUT[2383] <= 2766;PLUT[2384] <= 2750;PLUT[2385] <= 2733;PLUT[2386] <= 2717;PLUT[2387] <= 2701;PLUT[2388] <= 2685;PLUT[2389] <= 2669;PLUT[2390] <= 2653;PLUT[2391] <= 2637;PLUT[2392] <= 2621;PLUT[2393] <= 2606;PLUT[2394] <= 2590;PLUT[2395] <= 2575;PLUT[2396] <= 2559;PLUT[2397] <= 2544;PLUT[2398] <= 2529;PLUT[2399] <= 2514;PLUT[2400] <= 2499;PLUT[2401] <= 2484;PLUT[2402] <= 2469;PLUT[2403] <= 2454;PLUT[2404] <= 2440;PLUT[2405] <= 2425;PLUT[2406] <= 2411;PLUT[2407] <= 2396;PLUT[2408] <= 2382;PLUT[2409] <= 2368;PLUT[2410] <= 2354;PLUT[2411] <= 2340;PLUT[2412] <= 2326;PLUT[2413] <= 2312;PLUT[2414] <= 2298;PLUT[2415] <= 2284;PLUT[2416] <= 2271;PLUT[2417] <= 2257;PLUT[2418] <= 2244;PLUT[2419] <= 2230;PLUT[2420] <= 2217;PLUT[2421] <= 2204;PLUT[2422] <= 2191;PLUT[2423] <= 2177;PLUT[2424] <= 2164;PLUT[2425] <= 2152;PLUT[2426] <= 2139;PLUT[2427] <= 2126;PLUT[2428] <= 2113;PLUT[2429] <= 2101;PLUT[2430] <= 2088;PLUT[2431] <= 2076;PLUT[2432] <= 2063;PLUT[2433] <= 2051;PLUT[2434] <= 2039;PLUT[2435] <= 2027;PLUT[2436] <= 2015;PLUT[2437] <= 2002;PLUT[2438] <= 1991;PLUT[2439] <= 1979;PLUT[2440] <= 1967;PLUT[2441] <= 1955;PLUT[2442] <= 1943;PLUT[2443] <= 1932;PLUT[2444] <= 1920;PLUT[2445] <= 1909;PLUT[2446] <= 1898;PLUT[2447] <= 1886;PLUT[2448] <= 1875;PLUT[2449] <= 1864;PLUT[2450] <= 1853;PLUT[2451] <= 1842;PLUT[2452] <= 1831;PLUT[2453] <= 1820;PLUT[2454] <= 1809;PLUT[2455] <= 1798;PLUT[2456] <= 1787;PLUT[2457] <= 1777;PLUT[2458] <= 1766;PLUT[2459] <= 1756;PLUT[2460] <= 1745;PLUT[2461] <= 1735;PLUT[2462] <= 1724;PLUT[2463] <= 1714;PLUT[2464] <= 1704;PLUT[2465] <= 1694;PLUT[2466] <= 1683;PLUT[2467] <= 1673;PLUT[2468] <= 1663;PLUT[2469] <= 1654;PLUT[2470] <= 1644;PLUT[2471] <= 1634;PLUT[2472] <= 1624;PLUT[2473] <= 1614;PLUT[2474] <= 1605;PLUT[2475] <= 1595;PLUT[2476] <= 1586;PLUT[2477] <= 1576;PLUT[2478] <= 1567;PLUT[2479] <= 1557;PLUT[2480] <= 1548;PLUT[2481] <= 1539;PLUT[2482] <= 1530;PLUT[2483] <= 1521;PLUT[2484] <= 1512;PLUT[2485] <= 1503;PLUT[2486] <= 1494;PLUT[2487] <= 1485;PLUT[2488] <= 1476;PLUT[2489] <= 1467;PLUT[2490] <= 1458;PLUT[2491] <= 1450;PLUT[2492] <= 1441;PLUT[2493] <= 1432;PLUT[2494] <= 1424;PLUT[2495] <= 1415;PLUT[2496] <= 1407;PLUT[2497] <= 1398;PLUT[2498] <= 1390;PLUT[2499] <= 1382;PLUT[2500] <= 1374;PLUT[2501] <= 1365;PLUT[2502] <= 1357;PLUT[2503] <= 1349;PLUT[2504] <= 1341;PLUT[2505] <= 1333;PLUT[2506] <= 1325;PLUT[2507] <= 1317;PLUT[2508] <= 1309;PLUT[2509] <= 1302;PLUT[2510] <= 1294;PLUT[2511] <= 1286;PLUT[2512] <= 1278;PLUT[2513] <= 1271;PLUT[2514] <= 1263;PLUT[2515] <= 1256;PLUT[2516] <= 1248;PLUT[2517] <= 1241;PLUT[2518] <= 1233;PLUT[2519] <= 1226;PLUT[2520] <= 1219;PLUT[2521] <= 1211;PLUT[2522] <= 1204;PLUT[2523] <= 1197;PLUT[2524] <= 1190;PLUT[2525] <= 1183;PLUT[2526] <= 1176;PLUT[2527] <= 1169;PLUT[2528] <= 1162;PLUT[2529] <= 1155;PLUT[2530] <= 1148;PLUT[2531] <= 1141;PLUT[2532] <= 1134;PLUT[2533] <= 1127;PLUT[2534] <= 1121;PLUT[2535] <= 1114;PLUT[2536] <= 1107;PLUT[2537] <= 1101;PLUT[2538] <= 1094;PLUT[2539] <= 1088;PLUT[2540] <= 1081;PLUT[2541] <= 1075;PLUT[2542] <= 1068;PLUT[2543] <= 1062;PLUT[2544] <= 1056;PLUT[2545] <= 1049;PLUT[2546] <= 1043;PLUT[2547] <= 1037;PLUT[2548] <= 1031;PLUT[2549] <= 1024;PLUT[2550] <= 1018;PLUT[2551] <= 1012;PLUT[2552] <= 1006;PLUT[2553] <= 1000;PLUT[2554] <= 994;PLUT[2555] <= 988;PLUT[2556] <= 982;PLUT[2557] <= 977;PLUT[2558] <= 971;PLUT[2559] <= 965;PLUT[2560] <= 959;PLUT[2561] <= 953;PLUT[2562] <= 948;PLUT[2563] <= 942;PLUT[2564] <= 936;PLUT[2565] <= 931;PLUT[2566] <= 925;PLUT[2567] <= 920;PLUT[2568] <= 914;PLUT[2569] <= 909;PLUT[2570] <= 903;PLUT[2571] <= 898;PLUT[2572] <= 893;PLUT[2573] <= 887;PLUT[2574] <= 882;PLUT[2575] <= 877;PLUT[2576] <= 872;PLUT[2577] <= 866;PLUT[2578] <= 861;PLUT[2579] <= 856;PLUT[2580] <= 851;PLUT[2581] <= 846;PLUT[2582] <= 841;PLUT[2583] <= 836;PLUT[2584] <= 831;PLUT[2585] <= 826;PLUT[2586] <= 821;PLUT[2587] <= 816;PLUT[2588] <= 811;PLUT[2589] <= 806;PLUT[2590] <= 802;PLUT[2591] <= 797;PLUT[2592] <= 792;PLUT[2593] <= 787;PLUT[2594] <= 783;PLUT[2595] <= 778;PLUT[2596] <= 773;PLUT[2597] <= 769;PLUT[2598] <= 764;PLUT[2599] <= 759;PLUT[2600] <= 755;PLUT[2601] <= 750;PLUT[2602] <= 746;PLUT[2603] <= 742;PLUT[2604] <= 737;PLUT[2605] <= 733;PLUT[2606] <= 728;PLUT[2607] <= 724;PLUT[2608] <= 720;PLUT[2609] <= 715;PLUT[2610] <= 711;PLUT[2611] <= 707;PLUT[2612] <= 703;PLUT[2613] <= 698;PLUT[2614] <= 694;PLUT[2615] <= 690;PLUT[2616] <= 686;PLUT[2617] <= 682;PLUT[2618] <= 678;PLUT[2619] <= 674;PLUT[2620] <= 670;PLUT[2621] <= 666;PLUT[2622] <= 662;PLUT[2623] <= 658;PLUT[2624] <= 654;PLUT[2625] <= 650;PLUT[2626] <= 646;PLUT[2627] <= 642;PLUT[2628] <= 638;PLUT[2629] <= 635;PLUT[2630] <= 631;PLUT[2631] <= 627;PLUT[2632] <= 623;PLUT[2633] <= 620;PLUT[2634] <= 616;PLUT[2635] <= 612;PLUT[2636] <= 609;PLUT[2637] <= 605;PLUT[2638] <= 601;PLUT[2639] <= 598;PLUT[2640] <= 594;PLUT[2641] <= 591;PLUT[2642] <= 587;PLUT[2643] <= 584;PLUT[2644] <= 580;PLUT[2645] <= 577;PLUT[2646] <= 573;PLUT[2647] <= 570;PLUT[2648] <= 566;PLUT[2649] <= 563;PLUT[2650] <= 560;PLUT[2651] <= 556;PLUT[2652] <= 553;PLUT[2653] <= 550;PLUT[2654] <= 546;PLUT[2655] <= 543;PLUT[2656] <= 540;PLUT[2657] <= 537;PLUT[2658] <= 533;PLUT[2659] <= 530;PLUT[2660] <= 527;PLUT[2661] <= 524;PLUT[2662] <= 521;PLUT[2663] <= 518;PLUT[2664] <= 515;PLUT[2665] <= 512;PLUT[2666] <= 509;PLUT[2667] <= 505;PLUT[2668] <= 502;PLUT[2669] <= 499;PLUT[2670] <= 496;PLUT[2671] <= 494;PLUT[2672] <= 491;PLUT[2673] <= 488;PLUT[2674] <= 485;PLUT[2675] <= 482;PLUT[2676] <= 479;PLUT[2677] <= 476;PLUT[2678] <= 473;PLUT[2679] <= 470;PLUT[2680] <= 468;PLUT[2681] <= 465;PLUT[2682] <= 462;PLUT[2683] <= 459;PLUT[2684] <= 457;PLUT[2685] <= 454;PLUT[2686] <= 451;PLUT[2687] <= 448;PLUT[2688] <= 446;PLUT[2689] <= 443;PLUT[2690] <= 440;PLUT[2691] <= 438;PLUT[2692] <= 435;PLUT[2693] <= 433;PLUT[2694] <= 430;PLUT[2695] <= 427;PLUT[2696] <= 425;PLUT[2697] <= 422;PLUT[2698] <= 420;PLUT[2699] <= 417;PLUT[2700] <= 415;PLUT[2701] <= 412;PLUT[2702] <= 410;PLUT[2703] <= 407;PLUT[2704] <= 405;PLUT[2705] <= 403;PLUT[2706] <= 400;PLUT[2707] <= 398;PLUT[2708] <= 395;PLUT[2709] <= 393;PLUT[2710] <= 391;PLUT[2711] <= 388;PLUT[2712] <= 386;PLUT[2713] <= 384;PLUT[2714] <= 381;PLUT[2715] <= 379;PLUT[2716] <= 377;PLUT[2717] <= 375;PLUT[2718] <= 372;PLUT[2719] <= 370;PLUT[2720] <= 368;PLUT[2721] <= 366;PLUT[2722] <= 364;PLUT[2723] <= 361;PLUT[2724] <= 359;PLUT[2725] <= 357;PLUT[2726] <= 355;PLUT[2727] <= 353;PLUT[2728] <= 351;PLUT[2729] <= 349;PLUT[2730] <= 347;PLUT[2731] <= 345;PLUT[2732] <= 342;PLUT[2733] <= 340;PLUT[2734] <= 338;PLUT[2735] <= 336;PLUT[2736] <= 334;PLUT[2737] <= 332;PLUT[2738] <= 330;PLUT[2739] <= 328;PLUT[2740] <= 326;PLUT[2741] <= 325;PLUT[2742] <= 323;PLUT[2743] <= 321;PLUT[2744] <= 319;PLUT[2745] <= 317;PLUT[2746] <= 315;PLUT[2747] <= 313;PLUT[2748] <= 311;PLUT[2749] <= 309;PLUT[2750] <= 307;PLUT[2751] <= 306;PLUT[2752] <= 304;PLUT[2753] <= 302;PLUT[2754] <= 300;PLUT[2755] <= 298;PLUT[2756] <= 297;PLUT[2757] <= 295;PLUT[2758] <= 293;PLUT[2759] <= 291;PLUT[2760] <= 290;PLUT[2761] <= 288;PLUT[2762] <= 286;PLUT[2763] <= 284;PLUT[2764] <= 283;PLUT[2765] <= 281;PLUT[2766] <= 279;PLUT[2767] <= 278;PLUT[2768] <= 276;PLUT[2769] <= 274;PLUT[2770] <= 273;PLUT[2771] <= 271;PLUT[2772] <= 269;PLUT[2773] <= 268;PLUT[2774] <= 266;PLUT[2775] <= 265;PLUT[2776] <= 263;PLUT[2777] <= 262;PLUT[2778] <= 260;PLUT[2779] <= 258;PLUT[2780] <= 257;PLUT[2781] <= 255;PLUT[2782] <= 254;PLUT[2783] <= 252;PLUT[2784] <= 251;PLUT[2785] <= 249;PLUT[2786] <= 248;PLUT[2787] <= 246;PLUT[2788] <= 245;PLUT[2789] <= 243;PLUT[2790] <= 242;PLUT[2791] <= 240;PLUT[2792] <= 239;PLUT[2793] <= 238;PLUT[2794] <= 236;PLUT[2795] <= 235;PLUT[2796] <= 233;PLUT[2797] <= 232;PLUT[2798] <= 231;PLUT[2799] <= 229;PLUT[2800] <= 228;PLUT[2801] <= 226;PLUT[2802] <= 225;PLUT[2803] <= 224;PLUT[2804] <= 222;PLUT[2805] <= 221;PLUT[2806] <= 220;PLUT[2807] <= 218;PLUT[2808] <= 217;PLUT[2809] <= 216;PLUT[2810] <= 215;PLUT[2811] <= 213;PLUT[2812] <= 212;PLUT[2813] <= 211;PLUT[2814] <= 210;PLUT[2815] <= 208;PLUT[2816] <= 207;PLUT[2817] <= 206;PLUT[2818] <= 205;PLUT[2819] <= 203;PLUT[2820] <= 202;PLUT[2821] <= 201;PLUT[2822] <= 200;PLUT[2823] <= 199;PLUT[2824] <= 197;PLUT[2825] <= 196;PLUT[2826] <= 195;PLUT[2827] <= 194;PLUT[2828] <= 193;PLUT[2829] <= 191;PLUT[2830] <= 190;PLUT[2831] <= 189;PLUT[2832] <= 188;PLUT[2833] <= 187;PLUT[2834] <= 186;PLUT[2835] <= 185;PLUT[2836] <= 184;PLUT[2837] <= 183;PLUT[2838] <= 181;PLUT[2839] <= 180;PLUT[2840] <= 179;PLUT[2841] <= 178;PLUT[2842] <= 177;PLUT[2843] <= 176;PLUT[2844] <= 175;PLUT[2845] <= 174;PLUT[2846] <= 173;PLUT[2847] <= 172;PLUT[2848] <= 171;PLUT[2849] <= 170;PLUT[2850] <= 169;PLUT[2851] <= 168;PLUT[2852] <= 167;PLUT[2853] <= 166;PLUT[2854] <= 165;PLUT[2855] <= 164;PLUT[2856] <= 163;PLUT[2857] <= 162;PLUT[2858] <= 161;PLUT[2859] <= 160;PLUT[2860] <= 159;PLUT[2861] <= 158;PLUT[2862] <= 157;PLUT[2863] <= 156;PLUT[2864] <= 155;PLUT[2865] <= 154;PLUT[2866] <= 153;PLUT[2867] <= 152;PLUT[2868] <= 152;PLUT[2869] <= 151;PLUT[2870] <= 150;PLUT[2871] <= 149;PLUT[2872] <= 148;PLUT[2873] <= 147;PLUT[2874] <= 146;PLUT[2875] <= 145;PLUT[2876] <= 144;PLUT[2877] <= 144;PLUT[2878] <= 143;PLUT[2879] <= 142;PLUT[2880] <= 141;PLUT[2881] <= 140;PLUT[2882] <= 139;PLUT[2883] <= 138;PLUT[2884] <= 138;PLUT[2885] <= 137;PLUT[2886] <= 136;PLUT[2887] <= 135;PLUT[2888] <= 134;PLUT[2889] <= 134;PLUT[2890] <= 133;PLUT[2891] <= 132;PLUT[2892] <= 131;PLUT[2893] <= 130;PLUT[2894] <= 130;PLUT[2895] <= 129;PLUT[2896] <= 128;PLUT[2897] <= 127;PLUT[2898] <= 127;PLUT[2899] <= 126;PLUT[2900] <= 125;PLUT[2901] <= 124;PLUT[2902] <= 124;PLUT[2903] <= 123;PLUT[2904] <= 122;PLUT[2905] <= 121;PLUT[2906] <= 121;PLUT[2907] <= 120;PLUT[2908] <= 119;PLUT[2909] <= 118;PLUT[2910] <= 118;PLUT[2911] <= 117;PLUT[2912] <= 116;PLUT[2913] <= 116;PLUT[2914] <= 115;PLUT[2915] <= 114;PLUT[2916] <= 114;PLUT[2917] <= 113;PLUT[2918] <= 112;PLUT[2919] <= 112;PLUT[2920] <= 111;PLUT[2921] <= 110;PLUT[2922] <= 110;PLUT[2923] <= 109;PLUT[2924] <= 108;PLUT[2925] <= 108;PLUT[2926] <= 107;PLUT[2927] <= 106;PLUT[2928] <= 106;PLUT[2929] <= 105;PLUT[2930] <= 104;PLUT[2931] <= 104;PLUT[2932] <= 103;PLUT[2933] <= 103;PLUT[2934] <= 102;PLUT[2935] <= 101;PLUT[2936] <= 101;PLUT[2937] <= 100;PLUT[2938] <= 100;PLUT[2939] <= 99;PLUT[2940] <= 98;PLUT[2941] <= 98;PLUT[2942] <= 97;PLUT[2943] <= 97;PLUT[2944] <= 96;PLUT[2945] <= 95;PLUT[2946] <= 95;PLUT[2947] <= 94;PLUT[2948] <= 94;PLUT[2949] <= 93;PLUT[2950] <= 93;PLUT[2951] <= 92;PLUT[2952] <= 91;PLUT[2953] <= 91;PLUT[2954] <= 90;PLUT[2955] <= 90;PLUT[2956] <= 89;PLUT[2957] <= 89;PLUT[2958] <= 88;PLUT[2959] <= 88;PLUT[2960] <= 87;PLUT[2961] <= 87;PLUT[2962] <= 86;PLUT[2963] <= 86;PLUT[2964] <= 85;PLUT[2965] <= 85;PLUT[2966] <= 84;PLUT[2967] <= 84;PLUT[2968] <= 83;PLUT[2969] <= 83;PLUT[2970] <= 82;PLUT[2971] <= 82;PLUT[2972] <= 81;PLUT[2973] <= 81;PLUT[2974] <= 80;PLUT[2975] <= 80;PLUT[2976] <= 79;PLUT[2977] <= 79;PLUT[2978] <= 78;PLUT[2979] <= 78;PLUT[2980] <= 77;PLUT[2981] <= 77;PLUT[2982] <= 76;PLUT[2983] <= 76;PLUT[2984] <= 75;PLUT[2985] <= 75;PLUT[2986] <= 75;PLUT[2987] <= 74;PLUT[2988] <= 74;PLUT[2989] <= 73;PLUT[2990] <= 73;PLUT[2991] <= 72;PLUT[2992] <= 72;PLUT[2993] <= 71;PLUT[2994] <= 71;PLUT[2995] <= 71;PLUT[2996] <= 70;PLUT[2997] <= 70;PLUT[2998] <= 69;PLUT[2999] <= 69;PLUT[3000] <= 69;PLUT[3001] <= 68;PLUT[3002] <= 68;PLUT[3003] <= 67;PLUT[3004] <= 67;PLUT[3005] <= 66;PLUT[3006] <= 66;PLUT[3007] <= 66;PLUT[3008] <= 65;PLUT[3009] <= 65;PLUT[3010] <= 65;PLUT[3011] <= 64;PLUT[3012] <= 64;PLUT[3013] <= 63;PLUT[3014] <= 63;PLUT[3015] <= 63;PLUT[3016] <= 62;PLUT[3017] <= 62;PLUT[3018] <= 61;PLUT[3019] <= 61;PLUT[3020] <= 61;PLUT[3021] <= 60;PLUT[3022] <= 60;PLUT[3023] <= 60;PLUT[3024] <= 59;PLUT[3025] <= 59;PLUT[3026] <= 59;PLUT[3027] <= 58;PLUT[3028] <= 58;PLUT[3029] <= 58;PLUT[3030] <= 57;PLUT[3031] <= 57;PLUT[3032] <= 57;PLUT[3033] <= 56;PLUT[3034] <= 56;PLUT[3035] <= 55;PLUT[3036] <= 55;PLUT[3037] <= 55;PLUT[3038] <= 54;PLUT[3039] <= 54;PLUT[3040] <= 54;PLUT[3041] <= 54;PLUT[3042] <= 53;PLUT[3043] <= 53;PLUT[3044] <= 53;PLUT[3045] <= 52;PLUT[3046] <= 52;PLUT[3047] <= 52;PLUT[3048] <= 51;PLUT[3049] <= 51;PLUT[3050] <= 51;PLUT[3051] <= 50;PLUT[3052] <= 50;PLUT[3053] <= 50;PLUT[3054] <= 49;PLUT[3055] <= 49;PLUT[3056] <= 49;PLUT[3057] <= 49;PLUT[3058] <= 48;PLUT[3059] <= 48;PLUT[3060] <= 48;PLUT[3061] <= 47;PLUT[3062] <= 47;PLUT[3063] <= 47;PLUT[3064] <= 47;PLUT[3065] <= 46;PLUT[3066] <= 46;PLUT[3067] <= 46;PLUT[3068] <= 45;PLUT[3069] <= 45;PLUT[3070] <= 45;PLUT[3071] <= 45;
      out_couter_update_valid <= 0;
      out_pd_valid <= 0;
      out_pd_data <= 0;
      out_counter_data_new <= 0;
      out_id_data_next <= 0;
    end else begin
      case(pre_state)
        S_IDLE: begin
          if(in_next_valid)begin
            if(in_next_counter < C_MAGIC_NUMBER)begin             //if counter value is a small number, counter should be line way adding
              out_counter_data_new <= in_next_counter + in_next_length;
              out_couter_update_valid <= 1;
              out_pd_valid <= 0;
              out_id_data_next <= in_next_id;
            end else if(in_next_counter < 20'b1000_0000_0000_0000_0000) begin    //if C_Data should be inited, 20bits = 1 + 19 bits
              out_counter_data_new <= 20'b1000_0000_0100_1110_0010;        //C|=90(b1000...),c&=(1000...),c+=1250
              out_couter_update_valid <= 1;
              out_pd_valid <= 0;
              out_id_data_next <= in_next_id;
            end else if(set_plut_down == 0) begin                    //counter value is large number 
              pd_data_tmp <= PLUT[in_next_counter[18:0]];///////qsy
              next_length_tmp <= in_next_length;
              out_id_data_next <= in_next_id;
              out_couter_update_valid <= 0;
              out_pd_valid <= 0;
              out_counter_data_new <= in_next_counter;
            end else begin
			  lookup_add_bram <= in_next_counter[18:0];
			  next_length_tmp <= in_next_length;
              out_id_data_next <= in_next_id;
              out_couter_update_valid <= 0;
              out_pd_valid <= 0;
              out_counter_data_new <= in_next_counter;
			end
          end else begin
            out_pd_valid <= 0;
            out_couter_update_valid <= 0;
          end
        end
        S_ADD: begin
          out_pd_valid <= 0;
          out_couter_update_valid <= 0;
        end
        S_INITIAL: begin
          out_pd_valid <= 0;
          out_couter_update_valid <= 0;
        end
        S_CALCMUL: begin
          out_pd_data <= pd_data_tmp * next_length_tmp;
          out_pd_valid <= 1;
          out_couter_update_valid <= 0;
        end
		S_ENABLE: begin
          //
        end
	    S_LOOKUP: begin
          //
        end
	    S_CALCMUL2: begin
          out_pd_data <= lookup_data_bram * next_length_tmp;
          out_pd_valid <= 1;
          out_couter_update_valid <= 0;
        end
        S_RESET: begin
          out_pd_valid <= 0;
          out_couter_update_valid <= 0;
        end
      endcase
    end
  end
  
endmodule
